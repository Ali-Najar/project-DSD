library verilog;
use verilog.vl_types.all;
entity tb_parking is
end tb_parking;
